<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-301.048,-54.5889,-208.266,-100.449</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>-280,-5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_SMALL_INVERTER</type>
<position>-273,-5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-285,-67</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>-296.5,-32</position>
<gparam>LABEL_TEXT 4)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>-285,-70</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-285,-72.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>-285,-75</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-285,-79</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>-285,-82</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-285,-84.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>-285,-87</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AM_MUX_16x1</type>
<position>-274,-48</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_10</ID>11 </input>
<input>
<ID>IN_11</ID>15 </input>
<input>
<ID>IN_12</ID>15 </input>
<input>
<ID>IN_13</ID>15 </input>
<input>
<ID>IN_14</ID>15 </input>
<input>
<ID>IN_15</ID>15 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>11 </input>
<input>
<ID>IN_4</ID>11 </input>
<input>
<ID>IN_5</ID>11 </input>
<input>
<ID>IN_6</ID>15 </input>
<input>
<ID>IN_7</ID>15 </input>
<input>
<ID>IN_8</ID>11 </input>
<input>
<ID>IN_9</ID>11 </input>
<output>
<ID>OUT</ID>10 </output>
<input>
<ID>SEL_0</ID>7 </input>
<input>
<ID>SEL_1</ID>6 </input>
<input>
<ID>SEL_2</ID>5 </input>
<input>
<ID>SEL_3</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_MUX_4x1</type>
<position>-276,-83</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>14 </input>
<output>
<ID>OUT</ID>43 </output>
<input>
<ID>SEL_0</ID>42 </input>
<input>
<ID>SEL_1</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>-260.5,48</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>-279,-35</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>-279,-32.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>-259,-77.5</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>-279.5,-30</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>-279,-37.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-276,-61.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>-272,-61.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>-332.5,-5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>31</ID>
<type>DE_TO</type>
<position>-324,-5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-262,-73</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>-270,-48</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>-276,-76</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>-272,-75.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_TOGGLE</type>
<position>-292,-55.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>-291.5,-45</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_MUX_4x1</type>
<position>-276,-71</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>3 </input>
<output>
<ID>OUT</ID>44 </output>
<input>
<ID>SEL_0</ID>39 </input>
<input>
<ID>SEL_1</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_MUX_2x1</type>
<position>-262,-77.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>37 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>-332.5,10</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>-324.5,10</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>-275.5,49</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>-332.5,5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>DE_TO</type>
<position>-325,5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>-275.5,47</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>-260,42.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>-260.5,36.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>DA_FROM</type>
<position>-275.5,43.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>-275.5,41.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>71</ID>
<type>DA_FROM</type>
<position>-275.5,37.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>-275.5,35.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_SMALL_INVERTER</type>
<position>-265.5,43.5</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_SMALL_INVERTER</type>
<position>-267.5,37.5</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>-332.5,0</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>-325,0.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>80</ID>
<type>AE_OR3</type>
<position>-246,42.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<input>
<ID>IN_2</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>-241,42.5</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>-263,16</position>
<gparam>LABEL_TEXT f(ABCD)= (0,1,2,3,4,5,12,13,14,15)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>-262,9</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>-279.5,10</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>-279.5,7.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND2</type>
<position>-262,3</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>-262,-3</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>-279.5,4</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>-279.5,1</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>-280,-2</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_SMALL_INVERTER</type>
<position>-271,4</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AE_OR3</type>
<position>-249.5,3</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<input>
<ID>IN_2</ID>67 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>-244.5,3</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AE_SMALL_INVERTER</type>
<position>-272.5,7.5</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_SMALL_INVERTER</type>
<position>-272.5,10</position>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AE_SMALL_INVERTER</type>
<position>-271,1</position>
<input>
<ID>IN_0</ID>77 </input>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>-295.5,-13</position>
<gparam>LABEL_TEXT 3)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_AND2</type>
<position>-260,-15.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>DA_FROM</type>
<position>-277.5,-12.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>-277.5,-17</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>-260,-22.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>-277.5,-21.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>-277.5,-23.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_SMALL_INVERTER</type>
<position>-269,-21.5</position>
<input>
<ID>IN_0</ID>79 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_SMALL_INVERTER</type>
<position>-270.5,-17</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_SMALL_INVERTER</type>
<position>-270.5,-12.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_SMALL_INVERTER</type>
<position>-268.5,-23.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>168</ID>
<type>AE_OR2</type>
<position>-250,-19.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>-246,-19.5</position>
<input>
<ID>N_in0</ID>94 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>-296,16.5</position>
<gparam>LABEL_TEXT 2)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-278,-5,-275,-5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268,-5,-268,-4</points>
<intersection>-5 2</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268,-4,-265,-4</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-271,-5,-268,-5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-268 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-279,-68,-279,-67</points>
<connection>
<GID>49</GID>
<name>IN_3</name></connection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-283,-67,-279,-67</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-279 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-275.5,-38.5,-275.5,-37.5</points>
<connection>
<GID>16</GID>
<name>SEL_3</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-277,-37.5,-275.5,-37.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-275.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-274.5,-38.5,-274.5,-35</points>
<connection>
<GID>16</GID>
<name>SEL_2</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-277,-35,-274.5,-35</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-273.5,-38.5,-273.5,-32.5</points>
<connection>
<GID>16</GID>
<name>SEL_1</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-277,-32.5,-273.5,-32.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-273.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-272.5,-38.5,-272.5,-30</points>
<connection>
<GID>16</GID>
<name>SEL_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-277.5,-30,-272.5,-30</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-272.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-283,-70,-279,-70</points>
<connection>
<GID>49</GID>
<name>IN_2</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-330.5,-5,-326,-5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-271,-48,-271,-48</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>33</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-280,-55.5,-280,-45.5</points>
<intersection>-55.5 6</intersection>
<intersection>-54.5 15</intersection>
<intersection>-52.5 13</intersection>
<intersection>-51.5 12</intersection>
<intersection>-50.5 11</intersection>
<intersection>-47.5 10</intersection>
<intersection>-46.5 9</intersection>
<intersection>-45.5 14</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-290,-55.5,-277,-55.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-280,-46.5,-277,-46.5</points>
<connection>
<GID>16</GID>
<name>IN_9</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-280,-47.5,-277,-47.5</points>
<connection>
<GID>16</GID>
<name>IN_8</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-280,-50.5,-277,-50.5</points>
<connection>
<GID>16</GID>
<name>IN_5</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-280,-51.5,-277,-51.5</points>
<connection>
<GID>16</GID>
<name>IN_4</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-280,-52.5,-277,-52.5</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-280,-45.5,-277,-45.5</points>
<connection>
<GID>16</GID>
<name>IN_10</name></connection>
<intersection>-280 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-280,-54.5,-277,-54.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-280 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-279,-72.5,-279,-72</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-283,-72.5,-279,-72.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-279 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-283,-75,-279,-75</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-279 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-279,-75,-279,-74</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-75 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-279,-80,-279,-79</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-283,-79,-279,-79</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-279 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-283,-45,-283,-40.5</points>
<intersection>-45 1</intersection>
<intersection>-40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-289.5,-45,-283,-45</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-283 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-283,-40.5,-277,-40.5</points>
<connection>
<GID>16</GID>
<name>IN_15</name></connection>
<intersection>-283 0</intersection>
<intersection>-277 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-277,-53.5,-277,-40.5</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<connection>
<GID>16</GID>
<name>IN_6</name></connection>
<connection>
<GID>16</GID>
<name>IN_7</name></connection>
<connection>
<GID>16</GID>
<name>IN_11</name></connection>
<connection>
<GID>16</GID>
<name>IN_12</name></connection>
<connection>
<GID>16</GID>
<name>IN_13</name></connection>
<connection>
<GID>16</GID>
<name>IN_14</name></connection>
<intersection>-40.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-283,-82,-279,-82</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<connection>
<GID>17</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-330.5,10,-326.5,10</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-273.5,49,-263.5,49</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-330.5,5,-327,5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-273.5,47,-263.5,47</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-273.5,43.5,-267.5,43.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-263.5,43.5,-263,43.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-279,-84.5,-279,-84</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-283,-84.5,-279,-84.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-279 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-283,-87,-279,-87</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-279 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-279,-87,-279,-86</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-87 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-273.5,41.5,-263,41.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-265.5,37.5,-263.5,37.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-273.5,35.5,-263.5,35.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-330.5,0.5,-327,0.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-330.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-330.5,0,-330.5,0.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>0.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-252.5,44.5,-252.5,48</points>
<intersection>44.5 1</intersection>
<intersection>48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-252.5,44.5,-249,44.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-252.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-257.5,48,-252.5,48</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-257,42.5,-249,42.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-252.5,36.5,-252.5,40.5</points>
<intersection>36.5 2</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-252.5,40.5,-249,40.5</points>
<connection>
<GID>80</GID>
<name>IN_2</name></connection>
<intersection>-252.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-257.5,36.5,-252.5,36.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>-252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-243,42.5,-242,42.5</points>
<connection>
<GID>82</GID>
<name>N_in0</name></connection>
<connection>
<GID>80</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-273.5,37.5,-269.5,37.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>76</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-260,-77.5,-260,-77.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<connection>
<GID>53</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-276,-66,-276,-63.5</points>
<connection>
<GID>49</GID>
<name>SEL_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-275,-66,-275,-64.5</points>
<connection>
<GID>49</GID>
<name>SEL_0</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-272,-64.5,-272,-63.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-275,-64.5,-272,-64.5</points>
<intersection>-275 0</intersection>
<intersection>-272 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-262,-75,-262,-75</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-276,-78,-276,-78</points>
<connection>
<GID>17</GID>
<name>SEL_1</name></connection>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-275,-78,-275,-77.5</points>
<connection>
<GID>17</GID>
<name>SEL_0</name></connection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-275,-77.5,-272,-77.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-275 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268.5,-83,-268.5,-76.5</points>
<intersection>-83 2</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268.5,-76.5,-264,-76.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-268.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-273,-83,-268.5,-83</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-268.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-268.5,-78.5,-268.5,-71</points>
<intersection>-78.5 1</intersection>
<intersection>-71 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-268.5,-78.5,-264,-78.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-268.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-273,-71,-268.5,-71</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>-268.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-277.5,4,-273,4</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-269,4,-265,4</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-256,5,-256,9</points>
<intersection>5 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-256,5,-252.5,5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-256 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-259,9,-256,9</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-256 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-259,3,-252.5,3</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<connection>
<GID>128</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-256,-3,-256,1</points>
<intersection>-3 2</intersection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-256,1,-252.5,1</points>
<connection>
<GID>136</GID>
<name>IN_2</name></connection>
<intersection>-256 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-259,-3,-256,-3</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>-256 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-246.5,3,-245.5,3</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<connection>
<GID>136</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-278,-2,-265,-2</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-277.5,10,-274.5,10</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-270.5,10,-265,10</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-277.5,7.5,-274.5,7.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-270.5,8,-265,8</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-270.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-270.5,7.5,-270.5,8</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>8 1</intersection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-277.5,1,-273,1</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-269,1,-266.5,1</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>-266.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-266.5,1,-266.5,2</points>
<intersection>1 1</intersection>
<intersection>2 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-266.5,2,-265,2</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>-266.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-275.5,-21.5,-271,-21.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-267,-21.5,-263,-21.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-275.5,-12.5,-272.5,-12.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-268.5,-12.5,-263,-12.5</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-263 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-263,-14.5,-263,-12.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-275.5,-17,-272.5,-17</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>154</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-268.5,-16.5,-263,-16.5</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>-268.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-268.5,-17,-268.5,-16.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>-16.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-275.5,-23.5,-270.5,-23.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-266.5,-23.5,-263,-23.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-247,-19.5,-247,-19.5</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-18.5,-255,-15.5</points>
<intersection>-18.5 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-255,-18.5,-253,-18.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-257,-15.5,-255,-15.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-255,-22.5,-255,-20.5</points>
<intersection>-22.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-255,-20.5,-253,-20.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>-255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-257,-22.5,-255,-22.5</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>-255 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 1>
<page 2>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 2>
<page 3>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 3>
<page 4>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 4>
<page 5>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 5>
<page 6>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 6>
<page 7>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 7>
<page 8>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 8>
<page 9>
<PageViewport>0,126.574,938.642,-337.379</PageViewport></page 9></circuit>